library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Collision is
    port(
        clock : in std_logic;
        reset : in std_logic
    );
end entity Collision;


architecture Collisioin_ARCH of Collision is
    
begin
    
end architecture Collisioin_ARCH;
