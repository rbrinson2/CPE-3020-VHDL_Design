library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MineSweep is
    port(
        clk : in std_logic;
        rst : in std_logic
    );
end entity MineSweep;

architecture MineSweep_ARCH of MineSweep is
    
begin
    

    
end architecture MineSweep_ARCH;
