
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Intro_tb is
    port (
        sw: out std_ulogic_vector(3 downto 1)
    );
end entity Intro_tb;

architecture Intro_ARCH of Intro_tb is
    
begin
    
    
    
end architecture Intro_ARCH;