library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pract is
    port(
        clock : in std_logic;
        reset : in std_logic
    );
end entity pract;

architecture pract_ARCH of pract is
    
begin
    
end architecture pract_ARCH;
