
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MoveDetect_TB is
    port(
        clock : in std_logic;
        reset : in std_logic
    );
end entity MoveDetect_TB;


architecture MoveDetect_TB_ARCH of MoveDetect_TB is
    
begin
    
end architecture MoveDetect_TB_ARCH;
