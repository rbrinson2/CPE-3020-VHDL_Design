

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Randomizer_TB is
    port(
        clock : in std_logic;
        reset : in std_logic
    );
end entity Randomizer_TB;

architecture Randomizer_TB_ARCH of Randomizer is
    
begin
    
end architecture Randomizer_TB_ARCH;
