library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package MineSweepPackage is
    constant BOMBBUSWIDTH   : integer := 16;
    
    
    constant TILEBUSWIDTH   : integer := 16;
    constant MOVEWIDTH      : integer := 16;
    
end package MineSweepPackage;
