library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MineSweep_TB is
end entity MineSweep_TB;

architecture MineSweep_TB_ARCH of MineSweep_TB is
    
begin
    
    
end architecture MineSweep_TB_ARCH;

