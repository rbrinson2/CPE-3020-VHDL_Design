

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TileDriver is
    port(
        clock : in std_logic;
        reset : in std_logic
    );
end entity TileDriver;

architecture TileDriver_ARCH of TileDriver is
    
begin
    
end architecture TileDriver_ARCH;
